// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// sonata package

package sonata_pkg;

  localparam int unsigned GPIO_NUM = 3;
  localparam int unsigned UART_NUM = 5;
  localparam int unsigned I2C_NUM  = 2;
  localparam int unsigned SPI_NUM  = 5;

  localparam int unsigned SPI_CS_NUM = 4;

endpackage : sonata_pkg
